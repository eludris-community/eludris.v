module eludris

// Message is a struct that contains message data.
[noinit]
pub struct Message {
pub:
	author  string
	content string
}
