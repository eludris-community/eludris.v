module eludris

pub fn hello() string {
	return 'Hello!'
}
